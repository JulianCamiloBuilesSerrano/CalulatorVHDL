 LIBRARY IEEE;

USE ieee.std_logic_1164.all;
-------------------------------------------------------
-- result_1 son las decenas
-- result_2 son las unidades
ENTITY decen_uni IS
	PORT(		num				:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
								
				result_1 				:	OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0);
				
				result_2 				:	OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0));
				
END ENTITY decen_uni;
ARCHITECTURE behaviour OF decen_uni IS
SIGNAL v	: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL vector : STD_LOGIC_VECTOR(9 DOWNTO 0);

BEGIN
	--decenas
	WITH num SELECT
				result_1 <=
				-----------00-------------
				"0000" WHEN "00000000",
				"0000" WHEN "00000001",
				"0000" WHEN "00000010",
				"0000" WHEN "00000011",
				"0000" WHEN "00000100",
				"0000" WHEN "00000101",
				"0000" WHEN "00000110",
				"0000" WHEN "00000111",
				"0000" WHEN "00001000",
				"0000" WHEN "00001001",
				-----------10-------------
				"0001" WHEN "00001010",
				"0001" WHEN "00001011",
				"0001" WHEN "00001100",
				"0001" WHEN "00001101",
				"0001" WHEN "00001110",
				"0001" WHEN "00001111",
				"0001" WHEN "00010000",
				"0001" WHEN "00010001",
				"0001" WHEN "00010010",
				"0001" WHEN "00010011",
				-----------20-------------
				"0010" WHEN "00010100",
				"0010" WHEN "00010101",
				"0010" WHEN "00010110",
				"0010" WHEN "00010111",
				"0010" WHEN "00011000",
				"0010"WHEN "00011001",
				"0010" WHEN "00011010",
				"0010" WHEN "00011011",
				"0010" WHEN "00011100",
				"0010" WHEN "00011101",
				-----------30-------------
				"0011" WHEN "00011110",
				"0011" WHEN "00011111",
				"0011" WHEN "00100000",
				"0011" WHEN "00100001",
				"0011" WHEN "00100010",
				"0011" WHEN "00100011",
				"0011" WHEN "00100100",
				"0011" WHEN "00100101",
				"0011" WHEN "00100110",
				"0011" WHEN "00100111",
				-----------40-------------
				"0100" WHEN "00101000",
				"0100" WHEN "00101001",
				"0100" WHEN "00101010",
				"0100" WHEN "00101011",
				"0100" WHEN "00101100",
				"0100" WHEN "00101101",
				"0100" WHEN "00101110",
				"0100" WHEN "00101111",
				"0100" WHEN "00110000",
				"0100" WHEN "00110001",
				-----------50-------------
				"0101" WHEN "00110010",
				"0101" WHEN "00110011",
				"0101" WHEN "00110100",
				"0101" WHEN "00110101",
				"0101" WHEN "00110110",
				"0101" WHEN "00110111",
				"0101" WHEN "00111000",
				"0101" WHEN "00111001",
				"0101" WHEN "00111010",
				"0101" WHEN "00111011",
				-----------60-------------
				"0110" WHEN "00111100",
				"0110" WHEN "00111101",
				"0110" WHEN "00111110",
				"0110" WHEN "00111111",
				"0110" WHEN "01000000",
				"0110" WHEN "01000001",
				"0110" WHEN "01000010",
				"0110" WHEN "01000011",
				"0110" WHEN "01000100",
				"0110" WHEN "01000101",
				-----------70-------------
				"0111" WHEN "01000110",
				"0111" WHEN "01000111",
				"0111" WHEN "01001000",
				"0111" WHEN "01001001",
				"0111" WHEN "01001010",
				"0111" WHEN "01001011",
				"0111" WHEN "01001100",
				"0111" WHEN "01001101",
				"0111" WHEN "01001110",
				"0111" WHEN "01001111",
				-----------80-------------
				"1000" WHEN "01010000",
				"1000" WHEN "01010001",
				"1111" WHEN OTHERS;
		--unidades
		WITH num SELECT
				result_2 <=
				-----------00-------------
				"0000" WHEN "00000000",
				"0001" WHEN "00000001",
				"0010" WHEN "00000010",
				"0011" WHEN "00000011",
				"0100" WHEN "00000100",
				"0101" WHEN "00000101",
				"0110" WHEN "00000110",
				"0111" WHEN "00000111",
				"1000" WHEN "00001000",
				"1001" WHEN "00001001",
				-----------10-------------
				"0000" WHEN "00001010",
				"0001" WHEN "00001011",
				"0010" WHEN "00001100",
				"0011" WHEN "00001101",
				"0100" WHEN "00001110",
				"0101" WHEN "00001111",
				"0110" WHEN "00010000",
				"0111" WHEN "00010001",
				"1000" WHEN "00010010",
				"1001" WHEN "00010011",
				-----------20-------------
				"0000" WHEN "00010100",
				"0001" WHEN "00010101",
				"0010" WHEN "00010110",
				"0011" WHEN "00010111",
				"0100" WHEN "00011000",
				"0101" WHEN "00011001",
				"0110" WHEN "00011010",
				"0111" WHEN "00011011",
				"1000" WHEN "00011100",
				"1001" WHEN "00011101",
				-----------30-------------
				"0011" WHEN "00011110",
				"0011" WHEN "00011111",
				"0011" WHEN "00100000",
				"0011" WHEN "00100001",
				"0011" WHEN "00100010",
				"0011" WHEN "00100011",
				"0011" WHEN "00100100",
				"0011" WHEN "00100101",
				"0011" WHEN "00100110",
				"0011" WHEN "00100111",
				-----------40-------------
				"0000" WHEN "00101000",
				"0001" WHEN "00101001",
				"0010" WHEN "00101010",
				"0011" WHEN "00101011",
				"0100" WHEN "00101100",
				"0101" WHEN "00101101",
				"0110" WHEN "00101110",
				"0111" WHEN "00101111",
				"1000" WHEN "00110000",
				"1001" WHEN "00110001",
				-----------50-------------
				"0000" WHEN "00110010",
				"0001" WHEN "00110011",
				"0010" WHEN "00110100",
				"0011" WHEN "00110101",
				"0100" WHEN "00110110",
				"0101" WHEN "00110111",
				"0110" WHEN "00111000",
				"0111" WHEN "00111001",
				"1000" WHEN "00111010",
				"1001" WHEN "00111011",
				-----------60-------------
				"0000" WHEN "00111100",
				"0001" WHEN "00111101",
				"0010" WHEN "00111110",
				"0011" WHEN "00111111",
				"0100" WHEN "01000000",
				"0101" WHEN "01000001",
				"0110" WHEN "01000010",
				"0111" WHEN "01000011",
				"1000" WHEN "01000100",
				"1001" WHEN "01000101",
				-----------70-------------
				"0000" WHEN "01000110",
				"0001" WHEN "01000111",
				"0010" WHEN "01001000",
				"0011" WHEN "01001001",
				"0100" WHEN "01001010",
				"0101" WHEN "01001011",
				"0110" WHEN "01001100",
				"0111" WHEN "01001101",
				"1000" WHEN "01001110",
				"1001" WHEN "01001111",
				-----------80-------------
				"0000" WHEN "01010000",
				"0001" WHEN "01010001",
				"1111" WHEN OTHERS;
					
END behaviour;